module adder(
output[31:0] s,
input[31:0] a,
input[31:0] b,
input cin);

wire c4, c8, c12, c16, c20, c24, c28;

wire[3:0] g3_0, g7_4, g11_8, g15_12, g19_16, g23_20, g27_24, g31_28;
wire[3:0] p3_0, p7_4, p11_8, p15_12, p19_16, p23_20, p27_24, p31_28;
wire G3_0, G7_4, G11_8, G15_12, G19_16, G23_20, G27_24, G31_28;
wire P3_0, P7_4, P11_8, P15_12, P19_16, P23_20, P27_24, P31_28;

adder4_g_p_G_P_signals claSignal3_0(.g(g3_0), .p(p3_0), .G(G3_0), .P(P3_0), .a(a[3:0]), .b(b[3:0]));
adder4_g_p_G_P_signals claSignal7_4(.g(g7_4), .p(p7_4), .G(G7_4), .P(P7_4), .a(a[7:4]), .b(b[7:4]));
adder4_g_p_G_P_signals claSignal11_8(.g(g11_8), .p(p11_8), .G(G11_8), .P(P11_8), .a(a[11:8]), .b(b[11:8]));
adder4_g_p_G_P_signals claSignal15_12(.g(g15_12), .p(p15_12), .G(G15_12), .P(P15_12), .a(a[15:12]), .b(b[15:12]));
adder4_g_p_G_P_signals claSignal9_16(.g(g19_16), .p(p19_16), .G(G19_16), .P(P19_16), .a(a[19:16]), .b(b[19:16]));
adder4_g_p_G_P_signals claSignal23_20(.g(g23_20), .p(p23_20), .G(G23_20), .P(P23_20), .a(a[23:20]), .b(b[23:20]));
adder4_g_p_G_P_signals claSigna27_24(.g(g27_24), .p(p27_24), .G(G27_24), .P(P27_24), .a(a[27:24]), .b(b[27:24]));
adder4_g_p_G_P_signals claSigna31_28(.g(g31_28), .p(p31_28), .G(G31_28), .P(P31_28), .a(a[31:28]), .b(b[31:28]));

// c4 = G3_0 + P3_0*c0
wire P3_0c0;
and and1(P3_0c0, P3_0, cin);
or or1(c4, G3_0, P3_0c0);

// c8 = G7_4 + P7_4*G3_0 + P7_4*P3_0*c0
wire P7_4G3_0, P7_4P3_0c0;
and and2(P7_4G3_0, P7_4, G3_0);
and and3(P7_4P3_0c0, P7_4, P3_0c0);
or or2(c8, G7_4, P7_4G3_0, P7_4P3_0c0);

// c12 = G11_8 + P11_8*G7_4 + P11_8*P7_4*G3_0 + P11_8*P7_4*P3_0*c0
wire P11_8G7_4, P11_8P7_4G3_0, P11_8P7_4P3_0c0;
and and4(P11_8G7_4, P11_8, G7_4);
and and5(P11_8P7_4G3_0, P11_8, P7_4G3_0);
and and6(P11_8P7_4P3_0c0, P11_8, P7_4P3_0c0);
or or3(c12, G11_8, P11_8G7_4, P11_8P7_4G3_0, P11_8P7_4P3_0c0);

// c16 = G15_12 + P15_12*G11_8 + P15_12*P11_8*G7_4 + P15_12*P11_8*P7_4*G3_0 + P15_12P11_8*P7_4*P3_0*c0
wire P15_12G11_8, P15_12P11_8G7_4, P15_12P11_8P7_4G3_0, P15_12P11_8P7_4P3_0c0;
and and7(P15_12G11_8, P15_12, G11_8);
and and8(P15_12P11_8G7_4, P15_12, P11_8G7_4);
and and9(P15_12P11_8P7_4G3_0, P15_12, P11_8P7_4G3_0);
and and10(P15_12P11_8P7_4P3_0c0, P15_12, P11_8P7_4P3_0c0);
or or4(c16, G15_12, P15_12G11_8, P15_12P11_8G7_4, P15_12P11_8P7_4G3_0, P15_12P11_8P7_4P3_0c0);

// c20 = G19_16 + P19_16G15_12 + P19_16P15_12*G11_8 + P19_16P15_12*P11_8*G7_4 + P19_16P15_12*P11_8*P7_4*G3_0 + P19_16P15_12P11_8*P7_4*P3_0*c0
wire P19_16G15_12, P19_16P15_12G11_8, P19_16P15_12P11_8G7_4, P19_16P15_12P11_8P7_4G3_0, P19_16P15_12P11_8P7_4P3_0c0;
and and11(P19_16G15_12, P19_16, G15_12);
and and12(P19_16P15_12G11_8, P19_16, P15_12G11_8);
and and13(P19_16P15_12P11_8G7_4, P19_16, P15_12P11_8G7_4);
and and14(P19_16P15_12P11_8P7_4G3_0, P19_16, P15_12P11_8P7_4G3_0);
and and15(P19_16P15_12P11_8P7_4P3_0c0, P19_16, P15_12P11_8P7_4P3_0c0);
or or5(c20, G19_16, P19_16G15_12, P19_16P15_12G11_8, P19_16P15_12P11_8G7_4, P19_16P15_12P11_8P7_4G3_0, P19_16P15_12P11_8P7_4P3_0c0);

// c24 = G23_20 + P23_20G19_16 + P23_20P19_16G15_12 + P23_20P19_16P15_12*G11_8 + P23_20P19_16P15_12*P11_8*G7_4 + P23_20P19_16P15_12*P11_8*P7_4*G3_0 + P23_20P19_16P15_12P11_8*P7_4*P3_0*c0
wire P23_20G19_16, P23_20P19_16G15_12, P23_20P19_16P15_12G11_8, P23_20P19_16P15_12P11_8G7_4, P23_20P19_16P15_12P11_8P7_4G3_0, P23_20P19_16P15_12P11_8P7_4P3_0c0;
and and16(P23_20G19_16, P23_20, G19_16);
and and17(P23_20P19_16G15_12, P23_20, P19_16G15_12);
and and18(P23_20P19_16P15_12G11_8, P23_20, P19_16P15_12G11_8);
and and19(P23_20P19_16P15_12P11_8G7_4, P23_20, P19_16P15_12P11_8G7_4);
and and20(P23_20P19_16P15_12P11_8P7_4G3_0, P23_20, P19_16P15_12P11_8P7_4G3_0);
and and21(P23_20P19_16P15_12P11_8P7_4P3_0c0, P23_20, P19_16P15_12P11_8P7_4P3_0c0);
or or6(c24, G23_20, P23_20G19_16, P23_20P19_16G15_12, P23_20P19_16P15_12G11_8, P23_20P19_16P15_12P11_8G7_4, P23_20P19_16P15_12P11_8P7_4G3_0, P23_20P19_16P15_12P11_8P7_4P3_0c0);

// c28 = G27_24 + P27_24G23_20 + P27_24P23_20G19_16 + P27_24P23_20P19_16G15_12 + P27_24P23_20P19_16P15_12*G11_8 + P27_24P23_20P19_16P15_12*P11_8*G7_4 + P27_24P23_20P19_16P15_12*P11_8*P7_4*G3_0 + P27_24P23_20P19_16P15_12P11_8*P7_4*P3_0*c0
wire P27_24G23_20, P27_24P23_20G19_16, P27_24P23_20P19_16G15_12, P27_24P23_20P19_16P15_12G11_8, P27_24P23_20P19_16P15_12P11_8G7_4, P27_24P23_20P19_16P15_12P11_8P7_4G3_0, P27_24P23_20P19_16P15_12P11_8P7_4P3_0c0;
and and22(P27_24G23_20, P27_24, G23_20);
and and23(P27_24P23_20G19_16, P27_24, P23_20G19_16);
and and24(P27_24P23_20P19_16G15_12, P27_24, P23_20P19_16G15_12);
and and25(P27_24P23_20P19_16P15_12G11_8, P27_24, P23_20P19_16P15_12G11_8);
and and26(P27_24P23_20P19_16P15_12P11_8G7_4, P27_24, P23_20P19_16P15_12P11_8G7_4);
and and27(P27_24P23_20P19_16P15_12P11_8P7_4G3_0, P27_24, P23_20P19_16P15_12P11_8P7_4G3_0);
and and28(P27_24P23_20P19_16P15_12P11_8P7_4P3_0c0, P27_24, P23_20P19_16P15_12P11_8P7_4P3_0c0);
or or7(c28, G27_24, P27_24G23_20, P27_24P23_20G19_16, P27_24P23_20P19_16G15_12, P27_24P23_20P19_16P15_12G11_8, P27_24P23_20P19_16P15_12P11_8G7_4, P27_24P23_20P19_16P15_12P11_8P7_4G3_0, P27_24P23_20P19_16P15_12P11_8P7_4P3_0c0);

adder4_cla adder3_0(.s(s[3:0]), .g(g3_0), .p(p3_0), .a(a[3:0]), .b(b[3:0]), .cin(cin));
adder4_cla adder7_4(.s(s[7:4]), .g(g7_4), .p(p7_4), .a(a[7:4]), .b(b[7:4]), .cin(c4));
adder4_cla adder11_8(.s(s[11:8]), .g(g11_8), .p(p11_8), .a(a[11:8]), .b(b[11:8]), .cin(c8));
adder4_cla adder15_12(.s(s[15:12]), .g(g15_12), .p(p15_12), .a(a[15:12]), .b(b[15:12]), .cin(c12));
adder4_cla adder19_16(.s(s[19:16]), .g(g19_16), .p(p19_16), .a(a[19:16]), .b(b[19:16]), .cin(c16));
adder4_cla adder23_20(.s(s[23:20]), .g(g23_20), .p(p23_20), .a(a[23:20]), .b(b[23:20]), .cin(c20));
adder4_cla adder27_24(.s(s[27:24]), .g(g27_24), .p(p27_24), .a(a[27:24]), .b(b[27:24]), .cin(c24));
adder4_cla adder31_28(.s(s[31:28]), .g(g31_28), .p(p31_28), .a(a[31:28]), .b(b[31:28]), .cin(c28));

endmodule